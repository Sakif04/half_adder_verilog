
module fulladd ();

    assign a=0;
    assign b=1;
    assign c=a+b;


initial begin
  
  $display("heLloo"," ",c);
end

endmodule